// first code

m
and(out,in1,in2);    //whatever written first is the input rest all output     

endmodule