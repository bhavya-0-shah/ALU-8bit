module Invertereightbit 
(
input [7:0]A,
output [7:0]Ac
);

assign Ac= ~A;



endmodule

