module 4isto1mux
(
   input in1,
   input in2,
   input in3,
   input in4,
   input [1:0]s,
   output o


);

endmodule